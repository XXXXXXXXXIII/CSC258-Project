module decoder(KEYBOARDBUTTON, PLUGBOARDCHANGED);

    input [4:0] KEYBOARDBUTTON;
    input [49:0] PLUGBOARDCHANGED;
    
    output [25:0] OUT;
    
    reg OUT;
    
    always @(*)
    begin
	
	5'd0: OUT = PLUGBOARDCHANGED;
	5'd1: OUT = PLUGBOARDCHANGED;
	5'd2: OUT = PLUGBOARDCHANGED;
	5'd3: OUT = PLUGBOARDCHANGED;
	5'd4: OUT = PLUGBOARDCHANGED;
	5'd5: OUT = PLUGBOARDCHANGED;
	5'd6: OUT = PLUGBOARDCHANGED;
	5'd7: OUT = PLUGBOARDCHANGED;
	5'd8: OUT = PLUGBOARDCHANGED;
	5'd9: OUT = CHANGETO;
	5'd10: OUT = CHANGETO;
	5'd11: OUT = CHANGETO;
	5'd12: OUT = CHANGETO;
	5'd13: OUT = CHANGETO;
	5'd14: OUT = CHANGETO;
	5'd15: OUT = CHANGETO;
	5'd16: OUT = CHANGETO;
	5'd17: OUT = CHANGETO;
	5'd18: OUT = CHANGETO;
	5'd19: OUT = CHANGETO;
	5'd20: OUT = CHANGETO;
	5'd21: OUT = CHANGETO;
	5'd22: OUT = CHANGETO;
	5'd23: OUT = CHANGETO;
	5'd24: OUT = CHANGETO;
	5'd25: OUT = CHANGETO;
	
	default: OUT=5'd0;
    end


endmodule